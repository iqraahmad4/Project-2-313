module part4(SW, HEX0);
	
	input [2:0]SW;
	output [0:6]HEX0;
	assign HEX0=SW;
endmodule